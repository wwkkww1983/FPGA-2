module vga_display(
    input              vga_clk,                  //VGA����ʱ��
    input              sys_rst_n,                //��λ�ź�
    input	   [ 2:0]  switch,
    input      [11:0]  pixel_xpos,               //���ص������
    input      [11:0]  pixel_ypos,               //���ص�������  
      
    output reg [23:0]  pixel_data                //���ص�����
    );    
    
parameter  H_DISP = 12'd640;                    //�ֱ��ʡ�����
parameter  V_DISP = 12'd480;                    //�ֱ��ʡ�����

//wire
wire  [1:0]  switch_wave;
wire         switch_model;

//assign
assign {switch_wave , switch_model} = switch;

//������ʾ��������
localparam POS_X_wave  = 10'd188;                    //�ַ�������ʼ�������
localparam POS_Y_wave  = 10'd100;                    //�ַ�������ʼ��������
localparam WIDTH_wave  = 10'd264;                     //�ַ�������
localparam HEIGHT_wave = 10'd88;                     //�ַ�����߶�

//ģʽ��ʾ��������
localparam POS_X_model  = 10'd110;                    //�ַ�������ʼ�������
localparam POS_Y_model  = 10'd300;                    //�ַ�������ʼ��������
localparam WIDTH_model  = 10'd176;                     //�ַ�������
localparam HEIGHT_model = 10'd44;                     //�ַ�����߶�

localparam WHITE  = 24'b1111_1111_1111_1111_1111_1111;     //RGB565 ��ɫ
localparam BLACK  = 24'b0000_0000_0000_0000_0000_0000;     //RGB565 ��ɫ
localparam RED    = 24'b1111_1111_0000_0000_0000_0000;     //RGB565 ��ɫ
localparam GREEN  = 24'b0000_0000_1111_1111_0000_0000;     //RGB565 ��ɫ
localparam BLUE   = 24'b0000_0000_0000_0000_1111_1111;     //RGB565 ��ɫ

    
//*****************************************************
//**                    main code
//*****************************************************
//���ݵ�ǰ���ص�����ָ����ǰ���ص���ɫ���ݣ�����Ļ����ʾ����
reg  [263:0] char[87:0];                        //������ʾ����
reg  [175:0] char_model[43:0];                        //ģʽ��ʾ����

always @(posedge vga_clk) begin  //0���Ҳ�  01 ���ǲ� 2����   3��ݲ�
	case(switch_wave)
	2'd0:
		begin	
			char[0] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
			char[1] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[2] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[3] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[4] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[5] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[6] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[7] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[8] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[9] <=  264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[10] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[11] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[12] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[13] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[14] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[15] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[16] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[17] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[18] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[19] <= 264'h000000000000000000000000000000000000000000000000000000003C00000000;
            char[20] <= 264'h000000000000000000000000000000000000000000000000000000007F00000000;
            char[21] <= 264'h000000000000000000000000000000000003800000000000000000007F80000000;
            char[22] <= 264'h00000000000000000000000000000000000FE00000000000000000007FC0000000;
            char[23] <= 264'h00000FC0000000000000000000000000001FF00000000000000000007FC0000000;
            char[24] <= 264'h00003FFFFFFFFFFFFC0000001FC03FE0001FF00000000003000000007FC0000000;
            char[25] <= 264'h00007FFFFFFFFFFFFF8000007FFFFFE0001FF0000000000FC00000007FC0000000;
            char[26] <= 264'h0000FFFFFFFFFFFFFFC00000FFFFFFF0001FF8000000001FF00000007FC0000000;
            char[27] <= 264'h0000FFFFFFFFFFFFFFC00001FFFFFFE0001FF8000000001FF80078007FC0000000;
            char[28] <= 264'h0001FFFFFFFFFFFFFF800001FFFFFFE0001FF8000000001FFC00FC1F7FF8000000;
            char[29] <= 264'h0001FFFE007FFFFFFF000001FFF81FE0001FF8000000001FFF00FFFFFFFFFFC000;
            char[30] <= 264'h0003FF80007FE00000000001FF001FC1F87FF8000000000FFF80FFFFFFFFFFE000;
            char[31] <= 264'h0003FC00007FE00000000001F0001FC7FFFFFFFFFF800007FFE07FFFFFFFFFF000;
            char[32] <= 264'h0001E000007FC0000000000000001FC7FFFFFFFFFFF00003FFF07FFFFFFFFFF000;
            char[33] <= 264'h00000000003FC0000000000000001FCFFFFFFFFFFFE00001FFF87FC03F83FFF000;
            char[34] <= 264'h00000000003FC0000000000000001F8FFFFFFFFFFFE000003FFC7F003F8003F000;
            char[35] <= 264'h00000000003FC0000000000000001F8FFC03FFFFFFC0000000007E003F8003F000;
            char[36] <= 264'h00000000003FC0000000000000003F8FC007E1FFFF80000000007E003F8003F000;
            char[37] <= 264'h00000000003FC000000000001FFFFF8E000FF003FF00000000007E003F8003F000;
            char[38] <= 264'h00000000003FC000000000003FFFFF80001FF8007C00078000003E003F8003F000;
            char[39] <= 264'h00000000003FE000000000003FFFFF00003FF80000000FF000003E003F8003F000;
            char[40] <= 264'h00000078003FE000000000003FFFFF00007FF00000000FFC00003E003F8003E000;
            char[41] <= 264'h000000FC003FE000000000003FE0FF0000FFE00000000FFF00003E003F8003E000;
            char[42] <= 264'h000001FE003FFFFE000000003F801E0001FF802000000FFFC0003E307FFF83E000;
            char[43] <= 264'h000001FE003FFFFFC00000003F00000003FF00F800000FFFE0007E7FFFFFC1C000;
            char[44] <= 264'h000001FF003FFFFFE00000003F00000007FC03F800000FFFF8007E7FFFFFE08000;
            char[45] <= 264'h000001FF003FFFFFE00000003F0000001FF807FC00000FFFFE007E7FFFFFE00000;
            char[46] <= 264'h000000FF003FFFFFC00000003F0000007FE00FFC000007FFFF007E7FE03FE00000;
            char[47] <= 264'h000000FF003FFFFF800000003F000001FF801FFC000003FFFFC07E7E001FE00000;
            char[48] <= 264'h000000FF003FE000000000007F000007FE003FFC000000FFFF807E3E001FE00000;
            char[49] <= 264'h000000FE003FE000000000007F801E07FE007FF80000001FF8007C3F001FC00000;
            char[50] <= 264'h000000FE003FC000000000007FFFFF8FFFF8FFE00000000000007C3F803FC00000;
            char[51] <= 264'h0000007E003FC000000000007FFFFFCFFFFFFF800000000000007C1FC03F800000;
            char[52] <= 264'h0000007E003FC000000000007FFFFFC7FFFFFE00000000000000FC07F07F800000;
            char[53] <= 264'h0000007E003FC000000000007FFFFFC7FF87FC00000000000000FC03F8FF000000;
            char[54] <= 264'h0000007E003FC000000000007E00FFC1C01FF0800000000000E0F801FFFE000000;
            char[55] <= 264'h0000007E003FC0000000000000003FC0003FE1E00000000003E1F8007FFE000000;
            char[56] <= 264'h0000007E003FC0000000000000003FC0007F83F0000000001FC1F8003FFC000000;
            char[57] <= 264'h0000007E007FC0000000000000003FC001FF03F8000000007FC3F0001FF8000000;
            char[58] <= 264'h0000007E007FE0000000000000003FC003FC01FC00000003FF83F0000FFE000000;
            char[59] <= 264'h0000007E007FE0000000000000007FC00FF801FE0000000FFF07F0000FFF000000;
            char[60] <= 264'h0000007F007FFC000000000000007F801FF000FF0000007FFE0FE0001FFFC00000;
            char[61] <= 264'h0000007FFFFFFFFFF800000000007F803FE0007F800001FFFC1FE0003FFFF00000;
            char[62] <= 264'h03FFFFFFFFFFFFFFFFFFF8000000FF80FF80003FC00003FFF81FC0007FFFFC0000;
            char[63] <= 264'h07FFFFFFFFFFFFFFFFFFF8000000FF01FF80007FE00003FFF03FC000FF7FFF8000;
            char[64] <= 264'h0FFFFFFFFFFFFFFFFFFFF8000000FF03FFE000FFE00003FFE0FF8003FE3FFFE000;
            char[65] <= 264'h0FFFFFFFFFFFFFFFFFFFF0000001FE03FFF001FFF00003FF81FF000FFC1FFFFE00;
            char[66] <= 264'h1FFFFFFFFFFFFFFFFFFFF0000003FE07FFFC0FF3F80003FE03FF003FF80FFFFFE0;
            char[67] <= 264'h1FFFFFF800007FFFFFFFE0030007FC07FFFFFFE0FC0001F807FE00FFF007FFFFFC;
            char[68] <= 264'h1FFFF000000001FFFFFFE003E00FFC07FFFFFFC07C00000007F80FFFE001FFFFF8;
            char[69] <= 264'h1FFE00000000001FFFFFC001FFFFF801C1FFFF801C00000001E01FFF8000FFFFF0;
            char[70] <= 264'h1FE0000000000003FFFFC000FFFFF000007FFF000000000000003FFF00007FFFF0;
            char[71] <= 264'h0F000000000000007FFF80003FFFE000001FFE000000000000001FFC00003FFFE0;
            char[72] <= 264'h00000000000000000FFF00001FFFC0000007F8000000000000000FF000000FFFC0;
            char[73] <= 264'h000000000000000001FE000007FF0000000000000000000000000780000007FF80;
            char[74] <= 264'h00000000000000000030000001FC0000000000000000000000000000000001FF00;
            char[75] <= 264'h00000000000000000000000000000000000000000000000000000000000000FC00;
            char[76] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[77] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[78] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[79] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[80] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[81] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[82] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[83] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[84] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[85] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[86] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[87] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
		end
    2'd1:
        begin
            char[0]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[1]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[2]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[3]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[4]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[5]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[6]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[7]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[8]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[9]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[10] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[11] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[12] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[13] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[14] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[15] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[16] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[17] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[18] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[19] <= 264'h000000000000000000000000000000000000000000000000000000003C00000000;
            char[20] <= 264'h0000000000000000000000000000000003F0000000000000000000007F00000000;
            char[21] <= 264'h000000000000000000000000000000000FF0000000000000000000007F80000000;
            char[22] <= 264'h000000000000000000000000000000001FF0000000000000000000007FC0000000;
            char[23] <= 264'h000038000000000000000000000000007FF0000000000000000000007FC0000000;
            char[24] <= 264'h0001FFC0000000000000000000000003FFF0000000000003000000007FC0000000;
            char[25] <= 264'h0003FFFFE0000000600000000000000FFFF078000000000FC00000007FC0000000;
            char[26] <= 264'h0007FFFFFFFFFFFFFC0000000000007FFFFFFE000000001FF00000007FC0000000;
            char[27] <= 264'h000FFFFFFFFFFFFFFE000000700007FFFFFFFE000000001FF80078007FC0000000;
            char[28] <= 264'h000FFFFFFFFFFFFFFE0000007FFFFFFFF9FFFE000000001FFC00FC1F7FF8000000;
            char[29] <= 264'h000FFFFFFFFFFFFFFE0000007FFFFFFFE07FFE000000001FFF00FFFFFFFFFFC000;
            char[30] <= 264'h000FFFFFFFFFFFFFFE0000003FFFFFFF803FFE000000000FFF80FFFFFFFFFFE000;
            char[31] <= 264'h000FFFFFFFFFFFFFFC0000003FFFFFFE003FF80000000007FFE07FFFFFFFFFF000;
            char[32] <= 264'h000FFFFE000000FFF80000001FFFFFF0003FF00000000003FFF07FFFFFFFFFF000;
            char[33] <= 264'h0003C000000000000000000007FFFF00003FC00000000001FFF87FC03F83FFF000;
            char[34] <= 264'h00000000000000000000000001FFC000007F8000000000003FFC7F003F8003F000;
            char[35] <= 264'h0000000000000000000000000000000000FF80018000000000007E003F8003F000;
            char[36] <= 264'h00000000000000000000000000003F8003FF000FE000000000007E003F8003F000;
            char[37] <= 264'h00000000000000000000000000007FFFFFFFFFFFF000000000007E003F8003F000;
            char[38] <= 264'h00000000000000000000000000007FFFFFFFFFFFF000078000003E003F8003F000;
            char[39] <= 264'h00000000000000000000000000007FFFFFFFFFFFF0000FF000003E003F8003F000;
            char[40] <= 264'h00000000000000000000000000007FFFFFFFFFFFF0000FFC00003E003F8003E000;
            char[41] <= 264'h00000000000000000000000000007F801FFF001FF0000FFF00003E003F8003E000;
            char[42] <= 264'h00000FF80000007FC000000000007F0007FE000FF0000FFFC0003E307FFF83E000;
            char[43] <= 264'h00003FFFFFFFFFFFE000000000007F0007FE000FF0000FFFE0007E7FFFFFC1C000;
            char[44] <= 264'h00007FFFFFFFFFFFF000000000007F0007FE000FF0000FFFF8007E7FFFFFE08000;
            char[45] <= 264'h00007FFFFFFFFFFFF000000000007F000FFF000FF0000FFFFE007E7FFFFFE00000;
            char[46] <= 264'h0000FFFFFFFFFFFFF000000000007FFFFFFFFFFFF00007FFFF007E7FE03FE00000;
            char[47] <= 264'h0000FFFFFFFFFFFFE000000000007FFFFFFFFFFFF00003FFFFC07E7E001FE00000;
            char[48] <= 264'h0000FFFFF800003FC000000000007FFFFFFFFFFFF00000FFFF807E3E001FE00000;
            char[49] <= 264'h0000FFE0000000000000000000007FFFFFFFFFFFF000001FF8007C3F001FC00000;
            char[50] <= 264'h00007C00000000000000000000007FC01FFF001FF000000000007C3F803FC00000;
            char[51] <= 264'h00000000000000000000000000007F0007FE000FF000000000007C1FC03F800000;
            char[52] <= 264'h0000000000000000000000000000FF0007FE000FF00000000000FC07F07F800000;
            char[53] <= 264'h0000000000000000000000000000FF0007FE000FF00000000000FC03F8FF000000;
            char[54] <= 264'h0000000000000000000000000000FFC07FFFC0FFF000000000E0F801FFFE000000;
            char[55] <= 264'h0000000000000000000000000001FFFFFFFFFFFFF000000003E1F8007FFE000000;
            char[56] <= 264'h0000000000000000000000000001FFFFFFFFFFFFF00000001FC1F8003FFC000000;
            char[57] <= 264'h0000000000000000000000000003FFFFFFFFFFFFF00000007FC3F0001FF8000000;
            char[58] <= 264'h0000000001C00000000000000007FFFFFFFFFFFFF0000003FF83F0000FFE000000;
            char[59] <= 264'h00FFFFFFFFFFFFFFC0000000000FFFF03FFFE0FFF000000FFF07F0000FFF000000;
            char[60] <= 264'h03FFFFFFFFFFFFFFFFFF8000001FFE0007FE001FF000007FFE0FE0001FFFC00000;
            char[61] <= 264'h07FFFFFFFFFFFFFFFFFFF800003FFC0007FE000FF00001FFFC1FE0003FFFF00000;
            char[62] <= 264'h0FFFFFFFFFFFFFFFFFFFFC0000FFF80007FC000FF00003FFF81FC0007FFFFC0000;
            char[63] <= 264'h1FFFFFFFFFFFFFFFFFFFFC0003FFF80007FC000FF00003FFF03FC000FF7FFF8000;
            char[64] <= 264'h1FFFFFFFFFFFFFFFFFFFF8000FFFF00007FC000FF00003FFE0FF8003FE3FFFE000;
            char[65] <= 264'h3FFFFFF01FFFFFFFFFFFF800FFFFE00007FC000FF80003FF81FF000FFC1FFFFE00;
            char[66] <= 264'h3FFFE0000000FFFFFFFFF007FFFFC00007FC000FF80003FE03FF003FF80FFFFFE0;
            char[67] <= 264'h3FFC0000000003FFFFFFE00FFFFF800007FC000FF80001F807FE00FFF007FFFFFC;
            char[68] <= 264'h3FE000000000001FFFFFE00FFFFF000007FC000FF800000007F80FFFE001FFFFF8;
            char[69] <= 264'h1F80000000000001FFFFC007FFFE000007FC000FF800000001E01FFF8000FFFFF0;
            char[70] <= 264'h00000000000000003FFF0007FFFC000007FC000FF800000000003FFF00007FFFF0;
            char[71] <= 264'h000000000000000007FE0001FFF0000003FC000FF800000000001FFC00003FFFE0;
            char[72] <= 264'h000000000000000000E000003F80000003FC000FF000000000000FF000000FFFC0;
            char[73] <= 264'h0000000000000000000000000000000003F80007F000000000000780000007FF80;
            char[74] <= 264'h0000000000000000000000000000000001E00007E000000000000000000001FF00;
            char[75] <= 264'h00000000000000000000000000000000000000000000000000000000000000FC00;
            char[76] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[77] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[78] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[79] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[80] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[81] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[82] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[83] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[84] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[85] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[86] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[87] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
        end
    2'd2:
        begin
            char[0]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[1]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[2]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[3]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[4]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[5]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[6]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[7]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[8]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[9]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[10] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[11] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[12] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[13] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[14] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[15] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[16] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[17] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[18] <= 264'h000000000000000000000000000000000000000000000000000000000000000000; 
            char[19] <= 264'h0000000001C0000000000000000000000000000000000000000000003C00000000;
            char[20] <= 264'h0000000007E0000000000000000000000000000000000000000000007F00000000;
            char[21] <= 264'h000000000FF8000000000000000000000000000000000000000000007F80000000;
            char[22] <= 264'h000000001FFF000000000000000000000000000060000000000000007FC0000000;
            char[23] <= 264'h000000001FFFC000000000000000000000000001F8000000000000007FC0000000;
            char[24] <= 264'h000000001FFFF800000000000080000000000007F8000003000000007FC0000000;
            char[25] <= 264'h000000001FFFFF800000000003FFFFFFFF00000FFC00000FC00000007FC0000000;
            char[26] <= 264'h000000001FFFFFE00000000007FFFFFFFFC0003FFC00001FF00000007FC0000000;
            char[27] <= 264'h0000000003FFFFC0000000001FFFFFFFFFC000FFF800001FF80078007FC0000000;
            char[28] <= 264'h00000000000FFE00000000001FFFFFFFFFC003FFF000001FFC00FC1F7FF8000000;
            char[29] <= 264'h0000000000000000000000001FFFFFFFFFC00FFFE000001FFF00FFFFFFFFFFC000;
            char[30] <= 264'h0000000000000000000000001FFFFFFFF0007FFF8000000FFF80FFFFFFFFFFE000;
            char[31] <= 264'h007C00000000000000001C00000FE03F8001FFFC00000007FFE07FFFFFFFFFF000;
            char[32] <= 264'h01FFFFFFFFFFFFFFFFFFF800000FE03F800FFFF000000003FFF07FFFFFFFFFF000;
            char[33] <= 264'h03FFFFFFFFFFFFFFFFFFF800000FE03F803FFF8000000001FFF87FC03F83FFF000;
            char[34] <= 264'h07FFFFFFFFFFFFFFFFFFF800000FC03F807FFE00000000003FFC7F003F8003F000;
            char[35] <= 264'h07FFFFFFFFFFFFFFFFFFF000000FC03F803FC0000000000000007E003F8003F000;
            char[36] <= 264'h0FFFFFFFFFFFFFFFFFFFF000000FC03F800000002000000000007E003F8003F000;
            char[37] <= 264'h0FFFFFE001FFFFFFFFFFE000000FE03F80000001F000000000007E003F8003F000;
            char[38] <= 264'h0FFFC00001FF000FFFFFC000000FE03F80000003F800078000003E003F8003F000;
            char[39] <= 264'h1FF0000001FF00007FFF8000000FE03F80000007F8000FF000003E003F8003F000;
            char[40] <= 264'h0F00000003FE000007FF8000C00FE03F8000000FFC000FFC00003E003F8003E000;
            char[41] <= 264'h0000000003FE0000007E0003FFFFFFFFFFE0001FF8000FFF00003E003F8003E000;
            char[42] <= 264'h0000000003FE000000000007FFFFFFFFFFF0007FF8000FFFC0003E307FFF83E000;
            char[43] <= 264'h0000000007FF00000000000FFFFFFFFFFFF000FFE0000FFFE0007E7FFFFFC1C000;
            char[44] <= 264'h0000000007FFFE000000001FFFFFFFFFFFF003FF80000FFFF8007E7FFFFFE08000;
            char[45] <= 264'h000000000FFFFFFFE000001FFFFFFFFFFFE00FFF00000FFFFE007E7FFFFFE00000;
            char[46] <= 264'h000000000FFFFFFFF000001FFF8FE03F80003FFC000007FFFF007E7FE03FE00000;
            char[47] <= 264'h000000001FFFFFFFF000000E000FE03F8000FFF001E003FFFFC07E7E001FE00000;
            char[48] <= 264'h000000001FFFFFFFF0000000000FE03F8003FFC003F000FFFF807E3E001FE00000;
            char[49] <= 264'h000000003FF000FFF0000000000FE03F800FFF0003F8001FF8007C3F001FC00000;
            char[50] <= 264'h000000007FE0007FF0000000000FE03F803FFC0007F8000000007C3F803FC00000;
            char[51] <= 264'h00000000FFC0003FE0000000001FC03F807FE0000FF8000000007C1FC03F800000;
            char[52] <= 264'h00000001FF80003FE0000000001FC03F803F00001FF800000000FC07F07F800000;
            char[53] <= 264'h00000003FF00001FE0000000001FC03F800000003FF000000000FC03F8FF000000;
            char[54] <= 264'h00000007FE00001FC0000000003FC03F800000007FE0000000E0F801FFFE000000;
            char[55] <= 264'h0000000FFE00003FC0000000003FC03F80000000FFC0000003E1F8007FFE000000;
            char[56] <= 264'h0000001FFC00003FC0000000003F803F80000001FF8000001FC1F8003FFC000000;
            char[57] <= 264'h0000007FF800003FC0000000007F803F80000007FF0000007FC3F0001FF8000000;
            char[58] <= 264'h000000FFF000003F8000000000FF803F8000000FFE000003FF83F0000FFE000000;
            char[59] <= 264'h000003FFE000003F8000000000FF003F8000003FFC00000FFF07F0000FFF000000;
            char[60] <= 264'h000007FFC000007F8000000001FF003F8000007FF800007FFE0FE0001FFFC00000;
            char[61] <= 264'h00001FFF0000007F0000000007FE003F800001FFE00001FFFC1FE0003FFFF00000;
            char[62] <= 264'h00007FFE0000007F000000000FFE003F800007FFC00003FFF81FC0007FFFFC0000;
            char[63] <= 264'h0001FFFC000000FF000000007FFC003FC0001FFF800003FFF03FC000FF7FFF8000;
            char[64] <= 264'h0007FFF8000001FE00000003FFF8003FC0007FFE000003FFE0FF8003FE3FFFE000;
            char[65] <= 264'h003FFFF0400003FE0000001FFFF0003FC003FFFC000003FF81FF000FFC1FFFFE00;
            char[66] <= 264'h00FFFFC0700007FC0000001FFFE0003FC03FFFF0000003FE03FF003FF80FFFFFE0;
            char[67] <= 264'h07FFFF807C001FFC0000001FFFC0003FC1FFFFE0000001F807FE00FFF007FFFFFC;
            char[68] <= 264'h1FFFFE003F00FFF80000000FFF00003FCFFFFF800000000007F80FFFE001FFFFF8;
            char[69] <= 264'h1FFFF8003FFFFFF000000003FC00003FCFFFFE000000000001E01FFF8000FFFFF0;
            char[70] <= 264'h07FFE0001FFFFFE0000000000000003F87FFF0000000000000003FFF00007FFFF0;
            char[71] <= 264'h03FF80000FFFFFC0000000000000003F007F00000000000000001FFC00003FFFE0;
            char[72] <= 264'h0078000007FFFF80000000000000000C000000000000000000000FF000000FFFC0;
            char[73] <= 264'h0000000001FFFF000000000000000000000000000000000000000780000007FF80;
            char[74] <= 264'h00000000003FF8000000000000000000000000000000000000000000000001FF00;
            char[75] <= 264'h00000000000000000000000000000000000000000000000000000000000000FC00;
            char[76] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[77] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[78] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[79] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[80] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[81] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[82] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[83] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[84] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[85] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[86] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[87] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
        end
    2'd3:
        begin
            char[0]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[1]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[2]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[3]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[4]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[5]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[6]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[7]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[8]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[9]  <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[10] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[11] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[12] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[13] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[14] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[15] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[16] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[17] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[18] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[19] <= 264'h000000000000000000000000000000000000000000000000000000003C00000000;
            char[20] <= 264'h000000000000000000000000000000000000000000000000000000007F00000000;
            char[21] <= 264'h00000000000000000000000000000001F000000000000000000000007F80000000;
            char[22] <= 264'h000001C0000000000000000000000003F800000000000000000000007FC0000000;
            char[23] <= 264'h000003E000F8000001C0000000000007FC00000000000000000000007FC0000000;
            char[24] <= 264'h000007E001FFFFFFFFF0000000000007FC00000000000003000000007FC0000000;
            char[25] <= 264'h00000FE001FFFFFFFFF8000000000007FE0000000000000FC00000007FC0000000;
            char[26] <= 264'h00001FE001FFFFFFFFF800000007E007FE0000000000001FF00000007FC0000000;
            char[27] <= 264'h00003FC000FFFFFFFFF800000007F007FE0000000000001FF80078007FC0000000;
            char[28] <= 264'h00007F8000FF80007FF800000007F807FEFFFF800000001FFC00FC1F7FF8000000;
            char[29] <= 264'h0001FF0000FF000007F800000007F803FFFFFFC00000001FFF00FFFFFFFFFFC000;
            char[30] <= 264'h0003FFFF00FE000007F000000007F803FFFFFFC00000000FFF80FFFFFFFFFFE000;
            char[31] <= 264'h0007FFFFE0FF000007F000000007F803FFFFFFC000000007FFE07FFFFFFFFFF000;
            char[32] <= 264'h001FFFFFF0FF00000FF000000007F803FFFFFF0000000003FFF07FFFFFFFFFF000;
            char[33] <= 264'h003FFFFFF0FFFFFFFFF000000007F803FE00000000000001FFF87FC03F83FFF000;
            char[34] <= 264'h00FFFE03E0FFFFFFFFF000000007F803FE000000000000003FFC7F003F8003F000;
            char[35] <= 264'h03FFC00000FFFFFFFFF000000003F803FE0000000000000000007E003F8003F000;
            char[36] <= 264'h0FFF800000FFFFFFFFF000000003F803FE0000000000000000007E003F8003F000;
            char[37] <= 264'h3FFE000000FE00FFFFF000000003F803FE0000000000000000007E003F8003F000;
            char[38] <= 264'h3FFC000000FE007E07E000000007F803FE0000000000078000003E003F8003F000;
            char[39] <= 264'h1FF80000007E007E000000000007FFFFFFFFFFFFC0000FF000003E003F8003F000;
            char[40] <= 264'h1FE3FFFF007E007E00000003FFFFFFFFFFFFFFFFFFFC0FFC00003E003F8003E000;
            char[41] <= 264'h0FC7FFFFC07E007E00000007FFFFFFFFFFFFFFFFFFFC0FFF00003E003F8003E000;
            char[42] <= 264'h000FFFFFC07E007E0000000FFFFFFFFFFFFFFFFFFFF80FFFC0003E307FFF83E000;
            char[43] <= 264'h000FFFFF807FFCFE0000001FFFFFFFC1FFFFFFFFFFF00FFFE0007E7FFFFFC1C000;
            char[44] <= 264'h000FBF80007FFFFFFFFFF81FFFFFC001F803FFFFFFF00FFFF8007E7FFFFFE08000;
            char[45] <= 264'h00003F80007FFFFFFFFFF81FFFF00001F8000FFFFFE00FFFFE007E7FFFFFE00000;
            char[46] <= 264'h00003F8000FFFFFFFFFFF03FFC080003F80000FFFFC007FFFF007E7FE03FE00000;
            char[47] <= 264'h00003F8000FFFFFFFFFFF03FC01F0003F8000E0FFF8003FFFFC07E7E001FE00000;
            char[48] <= 264'h00003F8000FFFFFFFFFFE00C001F8003F8000F80FE0000FFFF807E3E001FE00000;
            char[49] <= 264'h00FFFFFE00FC007E03FFC000003F8007FC000FC00000001FF8007C3F001FC00000;
            char[50] <= 264'h01FFFFFFE0FC007E001F8000003FC007FC000FC00000000000007C3F803FC00000;
            char[51] <= 264'h03FFFFFFF0FC007E00060000001F800FFE000FE00000000000007C1FC03F800000;
            char[52] <= 264'h07FFFFFFF1FC007E00000000001F800FFF000FE0000000000000FC07F07F800000;
            char[53] <= 264'h07FFFF9FC1F8007E00000000001F801FFFC00FE0000000000000FC03F8FF000000;
            char[54] <= 264'h03803F8001F9E07E03F00000001F801FFFE00FC00000000000E0F801FFFE000000;
            char[55] <= 264'h00003F8001FBFFFFFFF80000001F803F9FF00FC00000000003E1F8007FFE000000;
            char[56] <= 264'h00003F8003FBFFFFFFFC0000001F807F8FF80FC0000000001FC1F8003FFC000000;
            char[57] <= 264'h00003F8003FFFFFFFFFC0000001F80FF03FC0FC0000000007FC3F0001FF8000000;
            char[58] <= 264'h00003F8047F7FFFFFFFC0000001F81FE01FE0FC000000003FF83F0000FFE000000;
            char[59] <= 264'h00003F83E7F7FC001FFC0000001F03FC007F0FC00000000FFF07F0000FFF000000;
            char[60] <= 264'h00003F8FCFF3F80003FC0000001F07F8003F8FC00000007FFE0FE0001FFFC00000;
            char[61] <= 264'h00003FFF8FF3F00001FC0000001F0FF0000FCFC0000001FFFC1FE0003FFFF00000;
            char[62] <= 264'h00007FFF1FE3F00001F80000001F3FC00007CFE0000003FFF81FC0007FFFFC0000;
            char[63] <= 264'h00007FFE3FE3F00001F80000003F3F000003CFE0000003FFF03FC000FF7FFF8000;
            char[64] <= 264'h00007FFC7FC3F00001F80000003F3C0000000FE0000003FFE0FF8003FE3FFFE000;
            char[65] <= 264'h00007FFCFF83F80001F80000003F000000001FE0000003FF81FF000FFC1FFFFE00;
            char[66] <= 264'h0000FFF9FF01F80001F80000007FFFFFFFFFFFE0000003FE03FF003FF80FFFFFE0;
            char[67] <= 264'h0000FFE1FE01F80003F80000007FFFFFFFFFFFF0000001F807FE00FFF007FFFFFC;
            char[68] <= 264'h0001FFC1F001FDFFFFF8000000FFFFFFFFFFFFF00000000007F80FFFE001FFFFF8;
            char[69] <= 264'h0000FF800001FFFFFFF8000000FFFFFFFFFFFFF00000000001E01FFF8000FFFFF0;
            char[70] <= 264'h0000FE000001FFFFFFF8000000FFFFFFFFFFFFF00000000000003FFF00007FFFF0;
            char[71] <= 264'h000078000001FFFFFFF8000000FFFFE0003FFFE00000000000001FFC00003FFFE0;
            char[72] <= 264'h000000000001FFFFFFF80000007FC000000007E00000000000000FF000000FFFC0;
            char[73] <= 264'h000000000000F8000FF00000001F0000000001800000000000000780000007FF80;
            char[74] <= 264'h000000000000C00001C0000000000000000000000000000000000000000001FF00;
            char[75] <= 264'h00000000000000000000000000000000000000000000000000000000000000FC00;
            char[76] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[77] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[78] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[79] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[80] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[81] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[82] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[83] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[84] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[85] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[86] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
            char[87] <= 264'h000000000000000000000000000000000000000000000000000000000000000000;
        end
    default:;
    endcase	
end

always @(posedge vga_clk) begin  //  0������  1��ɨƵ
    case(switch_model)
    1'b0:
        begin
            char_model[0]  <=176'h00000000000000000000000000000000000000000000;
            char_model[1]  <=176'h00000000000000000000000000000000000000000000;
            char_model[2]  <=176'h00000000000000000000000000000000000000000000;
            char_model[3]  <=176'h00000000000000000000000000000000000000000000;
            char_model[4]  <=176'h00000000000000000000000000000000000000000000;
            char_model[5]  <=176'h00000000000000000000000000000000000000000000;
            char_model[6]  <=176'h00000000000000000000000000000000000000000000;
            char_model[7]  <=176'h00000000000000000000000000000000000000000000;
            char_model[8]  <=176'h00000000000000000000000000000000000000000000;
            char_model[9]  <=176'h00000000000000000000000000000000000000000000;
            char_model[10] <=176'h0000000000000001E000000030000000000000380C00;
            char_model[11] <=176'h00000000000000F1F0F00000380387000000003C1E00;
            char_model[12] <=176'h007FFFFFF00000F1F0F00000780387000000003C1E00;
            char_model[13] <=176'h00FFFFFFF80000F1F1F00000781B87000000003C3E00;
            char_model[14] <=176'h01FFFFFFF8000071F1C00000783FFFFC0000003C3000;
            char_model[15] <=176'h01F0078000002001F000E006787FDFFC0000003C0000;
            char_model[16] <=176'h0080078000007FFFFFFFF00FFF838700001C1FFF0000;
            char_model[17] <=176'h000007800000FFFFFFFFF01FFF9FFFF0007FFFFFFF80;
            char_model[18] <=176'h000007800000F8000000F008781FFFF000FFFFFFFF80;
            char_model[19] <=176'h000007800000F07FFF8070007C1C00F000FFE03C0000;
            char_model[20] <=176'h000E07800000E07FFFC03000FE1FFFE000E0003C0000;
            char_model[21] <=176'h000F07FF8000E07803C03001FE1FFFE00000003E0000;
            char_model[22] <=176'h000F07FF8000E07801C03001FF1C00E00000001E0000;
            char_model[23] <=176'h000F07FF8000607FFFC03003BB9DFDE00019FF9F0000;
            char_model[24] <=176'h000F07800000403FFFC00007B8DFFFE0003FFFDF0000;
            char_model[25] <=176'h000F078000000001E000001F380E73C0007FFFCF8000;
            char_model[26] <=176'h000F0780000001FFFFFC003E380070000079F80F8000;
            char_model[27] <=176'h000F0780000001FFFFFC007E38FFFFFFE000F00FC000;
            char_model[28] <=176'h000F0780000001FFFFFC007C39FFFFFFE000F007E000;
            char_model[29] <=176'h000F0780000001C1E03C000039F8E0FFC000F003F000;
            char_model[30] <=176'h000F9FFC000001C1E03C00003980E20F8000FFFBFC00;
            char_model[31] <=176'h1FFFFFFFFFE003C1E03C00003801C7800000FFF9FF80;
            char_model[32] <=176'h3FFFFFFFFFC00381E03C00003803C7C000FFFFC0FFFE;
            char_model[33] <=176'h3FFFC3FFFFC00381E03C0000380F83F001FFFC007FFE;
            char_model[34] <=176'h7F80000FFF800781E03C0000387F00F801FF80001FFC;
            char_model[35] <=176'h38000000FF800F01E03C000038FE007C03F800000FF8;
            char_model[36] <=176'h000000001F000400E03C00003038000E0180000003F0;
            char_model[37] <=176'h000000000000000000000000000000000000000000C0;
            char_model[38] <=176'h00000000000000000000000000000000000000000000;
            char_model[39] <=176'h00000000000000000000000000000000000000000000;
            char_model[40] <=176'h00000000000000000000000000000000000000000000;
            char_model[41] <=176'h00000000000000000000000000000000000000000000;
            char_model[42] <=176'h00000000000000000000000000000000000000000000;
            char_model[43] <=176'h00000000000000000000000000000000000000000000;
        end
    1'b1:
        begin
            char_model[0]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[1]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[2]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[3]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[4]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[5]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[6]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[7]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[8]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[9]  <= 176'h00000000000000000000000000000000000000000000;
            char_model[10] <= 176'h003E0000000000000000000030000000000000380C00;
            char_model[11] <= 176'h003F0000000000E000000000380387000000003C1E00;
            char_model[12] <= 176'h003F0000000000F03FFFFE00780387000000003C1E00;
            char_model[13] <= 176'h003F00001E0038F07FFFFC00781B87000000003C3E00;
            char_model[14] <= 176'h003F0781FF003CFFF073FC00783FFFFC0000003C3000;
            char_model[15] <= 176'h063F0FFFFF803CFF80703806787FDFFC0000003C0000;
            char_model[16] <= 176'h0FFFFFFFFF801CF70870000FFF838700001C1FFF0000;
            char_model[17] <= 176'h1FFFFFFFFF8018F03FFFC01FFF9FFFF0007FFFFFFF80;
            char_model[18] <= 176'h1FFF1C003F8018F03FFFC008781FFFF000FFFFFFFF80;
            char_model[19] <= 176'h0C3F00003F01FFFFBE03C0007C1C00F000FFE03C0000;
            char_model[20] <= 176'h003F00003F03FFFFBCC1C000FE1FFFE000E0003C0000;
            char_model[21] <= 176'h003FF0003F03FFFF38E1C001FE1FFFE00000003E0000;
            char_model[22] <= 176'h007FFFFFFF0301E038E1C001FF1C00E00000001E0000;
            char_model[23] <= 176'h07FFFFFFFF0019E338E1C003BB9DFDE00019FF9F0000;
            char_model[24] <= 176'h1FFF1FFFFF0039E738E1C007B8DFFFE0003FFFDF0000;
            char_model[25] <= 176'h1FFE1FC03F0038EF38E1C01F380E73C0007FFFCF8000;
            char_model[26] <= 176'h1FFE00003F0070FE38E1C03E380070000079F80F8000;
            char_model[27] <= 176'h0E3E00003F00E0FC38E1C07E38FFFFFFE000F00FC000;
            char_model[28] <= 176'h003E00003F00C0F839C1C07C39FFFFFFE000F007E000;
            char_model[29] <= 176'h003E00003F0001F039C1C00039F8E0FFC000F003F000;
            char_model[30] <= 176'h003E0FFFFF8007E033D9C0003980E20F8000FFFBFC00;
            char_model[31] <= 176'h003F1FFFFF801FC007BE00003801C7800000FFF9FF80;
            char_model[32] <= 176'h003E3FFFFF807F000F3F00003803C7C000FFFFC0FFFE;
            char_model[33] <= 176'hF87E3FFFFF03FE003E1F8000380F83F001FFFC007FFE;
            char_model[34] <= 176'h7FFE18000003F807FC07C000387F00F801FF80001FFC;
            char_model[35] <= 176'h3FFC00000001E007F803E00038FE007C03F800000FF8;
            char_model[36] <= 176'h1FF8000000000003E000F0003038000E0180000003F0;
            char_model[37] <= 176'h03E000000000000000001000000000000000000000C0;
            char_model[38] <= 176'h00000000000000000000000000000000000000000000;
            char_model[39] <= 176'h00000000000000000000000000000000000000000000;
            char_model[40] <= 176'h00000000000000000000000000000000000000000000;
            char_model[41] <= 176'h00000000000000000000000000000000000000000000;
            char_model[42] <= 176'h00000000000000000000000000000000000000000000;
            char_model[43] <= 176'h00000000000000000000000000000000000000000000;
        end
    default:;
    endcase
end
//wire define   
wire [ 9:0] x_cnt_wave;
wire [ 9:0] y_cnt_wave;
wire [11:0] x_cnt_model;
wire [11:0] y_cnt_model;

assign x_cnt_wave  = pixel_xpos - POS_X_wave;              //���ص�����ڲ�����ʾ������ʼ��ˮƽ����
assign y_cnt_wave  = pixel_ypos - POS_Y_wave;              //���ص�����ڲ�����ʾ������ʼ����ֱ����
assign x_cnt_model = pixel_xpos - POS_X_model;              //���ص������ģʽ��ʾ������ʼ��ˮƽ����
assign y_cnt_model = pixel_ypos - POS_Y_model;              //���ص������ģʽ��ʾ������ʼ����ֱ����

always @(posedge vga_clk or negedge sys_rst_n) begin        //��ʾ
    if (!sys_rst_n) 
        pixel_data <= BLACK;
    else if((pixel_xpos >= POS_X_wave) && (pixel_xpos < POS_X_wave + WIDTH_wave)
          && (pixel_ypos >= POS_Y_wave) && (pixel_ypos < POS_Y_wave + HEIGHT_wave)) 
        begin
            if(char[y_cnt_wave][10'd263 - x_cnt_wave])
                pixel_data <= WHITE;              //�����ַ�Ϊ��ɫ
            else
                pixel_data <= BLACK;             //�����ַ����򱳾�Ϊ��ɫ      
        end
    else if((pixel_xpos >= POS_X_model) && (pixel_xpos < POS_X_model + WIDTH_model)
          && (pixel_ypos >= POS_Y_model) && (pixel_ypos < POS_Y_model + HEIGHT_model))
        begin
            if(char_model[y_cnt_model][10'd175 - x_cnt_model])
                pixel_data <= WHITE;              //�����ַ�Ϊ��ɫ
            else
                pixel_data <= BLACK;             //�����ַ����򱳾�Ϊ��ɫ      
        end
    else
            pixel_data <= BLACK;                //������Ļ����Ϊ��ɫ
end


endmodule 